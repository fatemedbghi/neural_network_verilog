`timescale 1ns / 1ns

module NeuraNetworkController();


endmodule
