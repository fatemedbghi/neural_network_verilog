`timescale 1ns / 1ns

module Neuron10 # (
		parameter DW = 8,
		parameter DW_VEC = 8,
		parameter O_VEC = 21)
		(input wire clk, rst, start, output wire [79:0] out);

		
		
endmodule
