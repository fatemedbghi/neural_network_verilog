`timescale 1ns / 1ps

module NeuralNetworkDataPath(input [61:0] test_data, output integer test_out);


endmodule
